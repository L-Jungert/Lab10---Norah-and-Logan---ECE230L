module demux2(
    input [1:0] data,
    input [1:0] sel,
    output reg [1:0] A,
    output reg [1:0] B, 
    output reg [1:0] C, 
    output reg [1:0] D
);
    always @(*) begin
        case (sel)
            2'b00: {D,C,B,A} <= {2'b0,2'b0,2'b0,data};
            2'b01: {D,C,B,A} <= {2'b0,2'b0,data,2'b0};
            2'b10: {D,C,B,A} <= {2'b0,data,2'b0,2'b0};
            2'b11: {D,C,B,A} <= {data,2'b0,2'b0,2'b0};
        endcase
    end
endmodule
